module SEXT(
    input wire [31:0] inst,
    input wire [2:0]  sext_op,
    output wire [31:0] ext
);

// 000 ---> no imm
// 001 ---> 0000_0000_0000_0000_0000_inst[31:20]
// 010 ---> 0000_0000_0000_0000_0000_inst[31:25|11:7]
// 011 ---> 0000_0000_0000_0000_000_inst[31|7|30:25|11:8]_0;
// 100 ---> inst[31:12]|0000_0000_0000;
// 101 ---> 0000_0000_000_inst[31|19:12|20|30|21]_0
assign ext = (sext_op == 3'b000) ? 32'b0 :
             (sext_op == 3'b001) ? (inst[31] == 1'b1 ? {20'b1111_1111_1111_1111_1111, inst[31:20]} : {20'b0000_0000_0000_0000_0000, inst[31:20]}) :
             (sext_op == 3'b010) ? (inst[31] == 1'b1 ? {20'b1111_1111_1111_1111_1111, inst[31:25], inst[11:7]} : {20'b0000_0000_0000_0000_0000, inst[31:25], inst[11:7]})   :
             (sext_op == 3'b011) ? (inst[31] == 1'b1 ? {19'b1111_1111_1111_1111_111, inst[31], inst[7], inst[30:25], inst[11:8], 1'b0} : {19'b0000_0000_0000_0000_000, inst[31], inst[7], inst[30:25], inst[11:8], 1'b0})  :
             (sext_op == 3'b100) ? {inst[31:12], 12'b0000_0000_0000} : 
                                   (inst[31] == 1'b1 ? {11'b1111_1111_111, inst[31], inst[19:12], inst[20], inst[30:21], 1'b0} : {11'b0000_0000_000, inst[31], inst[19:12], inst[20], inst[30:21], 1'b0});
endmodule